module Main(input );

