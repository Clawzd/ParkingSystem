module Main(input normal_spaces);

  wire D1= normal_spaces / 10 ;
  wire D0= normal_spaces % 10 ;
