module Main(input [4:0]normal_spaces);

  wire [3:0]D1= normal_spaces/10 ;
  wire [3:0]D0= normal_spaces%10 ;
