module Main(input clk, n_entry, n_exit, h_entry , h_exit , reset, output );

